`default_nettype none

module shifter #(
   parameter N=32
)(
   input  wire signed [N-1:0] IN,
   input  wire        [$clog2(N)-1:0] shamt, // arredondando para log2
   input  wire left, logical,
   output wire [N-1:0] OUT
);

   assign OUT = left ?  (IN << shamt) :
                        (logical ? IN >> shamt : IN >>> shamt);

endmodule